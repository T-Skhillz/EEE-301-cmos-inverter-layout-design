magic
tech sky130A
magscale 1 2
timestamp 1770660156
<< metal1 >>
rect -2994 3202 -838 3206
rect -2994 3198 -626 3202
rect -502 3198 598 3206
rect -2994 2790 598 3198
rect -1404 2194 -998 2790
rect -2266 2102 -2122 2120
rect -2266 2047 -2247 2102
rect -2159 2047 -2122 2102
rect -2266 2032 -2122 2047
rect -2000 2036 -1800 2052
rect -2000 1944 -1980 2036
rect -1820 1944 -1800 2036
rect -2000 1932 -1800 1944
rect -2302 1420 -2102 1474
rect -2660 1380 -1260 1420
rect -2660 1300 -2620 1380
rect -2500 1320 -1420 1380
rect -1340 1320 -1260 1380
rect -2500 1300 -1260 1320
rect -2660 1280 -1260 1300
rect -2302 1274 -2102 1280
rect -1264 947 -1149 982
rect -1698 700 -1498 900
rect -1360 860 -1240 880
rect -820 860 -720 862
rect -1360 760 -1340 860
rect -1260 760 -1240 860
rect -1360 720 -1240 760
rect -1108 759 -720 860
rect -820 216 -720 759
rect -3002 -200 590 216
<< via1 >>
rect -2247 2047 -2159 2102
rect -1980 1944 -1820 2036
rect -2620 1300 -2500 1380
rect -1420 1320 -1340 1380
rect -1340 760 -1260 860
<< metal2 >>
rect -2624 2122 -2481 2123
rect -2624 2120 -2353 2122
rect -2624 2102 -2122 2120
rect -2624 2047 -2247 2102
rect -2159 2047 -2122 2102
rect -2624 2034 -2122 2047
rect -2624 2032 -2481 2034
rect -2368 2032 -2122 2034
rect -2000 2036 -1800 2052
rect -2620 1420 -2500 2032
rect -2000 1944 -1980 2036
rect -1820 1944 -1800 2036
rect -2660 1380 -2460 1420
rect -2660 1300 -2620 1380
rect -2500 1300 -2460 1380
rect -2660 1280 -2460 1300
rect -2620 1120 -2500 1280
rect -2000 900 -1800 1944
rect -1260 1283 -1100 1420
rect -1264 1280 -1100 1283
rect -1264 947 -1159 1280
rect -2000 880 -1281 900
rect -2000 860 -1240 880
rect -2000 760 -1340 860
rect -1260 760 -1240 860
rect -2000 720 -1240 760
rect -2000 700 -1281 720
rect -2000 698 -1800 700
<< rmetal2 >>
rect -1740 1380 -1260 1420
rect -1740 1320 -1420 1380
rect -1340 1320 -1260 1380
rect -1740 1283 -1260 1320
rect -1740 1280 -1264 1283
use sky130_fd_pr__nfet_01v8_66VXEL  sky130_fd_pr__nfet_01v8_66VXEL_0
timestamp 1770646034
transform 1 0 -1200 0 1 810
box -276 -310 276 310
use sky130_fd_pr__pfet_01v8_89MGVZ  sky130_fd_pr__pfet_01v8_89MGVZ_0
timestamp 1770646034
transform 0 1 -1185 -1 0 2070
box -276 -1219 276 1219
<< labels >>
flabel metal1 -1300 2904 -1100 3104 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 -1296 -112 -1096 88 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 -2302 1274 -2102 1474 0 FreeSans 256 0 0 0 Vin
port 0 nsew
flabel metal1 -1698 700 -1498 900 0 FreeSans 256 0 0 0 Vout
port 2 nsew
<< end >>
